module NOC #(parameter flit_width=16,MAX_Packet_NUM=8,Flit_size = 16, REQ_size = 3,NUM_OF_ROUTERS = 9)
(
input    wire                                               clk,                                                                            
input    wire                                               rst,
//PE ports
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_VALID_i,
input    wire   [NUM_OF_ROUTERS*flit_width-1:0]             PE_FLIT_i,
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_VC_0_RESERVED_i,
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_VC_1_RESERVED_i,
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_VC_2_RESERVED_i,
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_VC_3_RESERVED_i,
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_ON_OFF_0_i,
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_ON_OFF_1_i,
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_ON_OFF_2_i,
input    wire   [NUM_OF_ROUTERS-1:0]                        PE_ON_OFF_3_i,
//north ports
input    wire   [(3*flit_width)-1:0]                        in_N_FLIT_i,
input    wire   [2:0]                                       in_N_VALID_i,        
input    wire   [2:0]                                       in_N_VC_0_RESERVED_i,
input    wire   [2:0]                                       in_N_VC_1_RESERVED_i,
input    wire   [2:0]                                       in_N_VC_2_RESERVED_i,
input    wire   [2:0]                                       in_N_VC_3_RESERVED_i,
input    wire   [2:0]                                       in_N_ON_OFF_0_i,
input    wire   [2:0]                                       in_N_ON_OFF_1_i,
input    wire   [2:0]                                       in_N_ON_OFF_2_i,
input    wire   [2:0]                                       in_N_ON_OFF_3_i,
//south ports													 
input    wire   [(3*flit_width)-1:0]                        in_S_FLIT_i,
input    wire   [2:0]                                       in_S_VALID_i,        
input    wire   [2:0]                                       in_S_VC_0_RESERVED_i,
input    wire   [2:0]                                       in_S_VC_1_RESERVED_i,
input    wire   [2:0]                                       in_S_VC_2_RESERVED_i,
input    wire   [2:0]                                       in_S_VC_3_RESERVED_i,
input    wire   [2:0]                                       in_S_ON_OFF_0_i,
input    wire   [2:0]                                       in_S_ON_OFF_1_i,
input    wire   [2:0]                                       in_S_ON_OFF_2_i,
input    wire   [2:0]                                       in_S_ON_OFF_3_i,
//weast ports													 
input    wire   [(3*flit_width)-1:0]                        in_W_FLIT_i,
input    wire   [2:0]                                       in_W_VALID_i,        
input    wire   [2:0]                                       in_W_VC_0_RESERVED_i,
input    wire   [2:0]                                       in_W_VC_1_RESERVED_i,
input    wire   [2:0]                                       in_W_VC_2_RESERVED_i,
input    wire   [2:0]                                       in_W_VC_3_RESERVED_i,
input    wire   [2:0]                                       in_W_ON_OFF_0_i,
input    wire   [2:0]                                       in_W_ON_OFF_1_i,
input    wire   [2:0]                                       in_W_ON_OFF_2_i,
input    wire   [2:0]                                       in_W_ON_OFF_3_i,
//east ports													 
input    wire   [(3*flit_width)-1:0]                        in_E_FLIT_i,
input    wire   [2:0]                                       in_E_VALID_i,        
input    wire   [2:0]                                       in_E_VC_0_RESERVED_i,
input    wire   [2:0]                                       in_E_VC_1_RESERVED_i,
input    wire   [2:0]                                       in_E_VC_2_RESERVED_i,
input    wire   [2:0]                                       in_E_VC_3_RESERVED_i,
input    wire   [2:0]                                       in_E_ON_OFF_0_i,
input    wire   [2:0]                                       in_E_ON_OFF_1_i,
input    wire   [2:0]                                       in_E_ON_OFF_2_i,
input    wire   [2:0]                                       in_E_ON_OFF_3_i,

//outputs 
//PE ports
output   wire   [NUM_OF_ROUTERS*flit_width-1:0]          PE_FLIT_o,               
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_VALID_O,
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_VC_0_RESERVED_O,
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_VC_1_RESERVED_O,
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_VC_2_RESERVED_O,
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_VC_3_RESERVED_O,
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_ON_OFF_0_O,
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_ON_OFF_1_O,
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_ON_OFF_2_O,
output   wire   [NUM_OF_ROUTERS-1:0]                     PE_ON_OFF_3_O,
//north ports
output   wire   [(3*flit_width)-1:0]                     out_N_FLIT_o,
output   wire   [2:0]                                    out_N_VALID_O,
output   wire   [2:0]                                    out_N_VC_0_RESERVED_O,
output   wire   [2:0]                                    out_N_VC_1_RESERVED_O,
output   wire   [2:0]                                    out_N_VC_2_RESERVED_O,
output   wire   [2:0]                                    out_N_VC_3_RESERVED_O,
output   wire   [2:0]                                    out_N_ON_OFF_0_O,
output   wire   [2:0]                                    out_N_ON_OFF_1_O,
output   wire   [2:0]                                    out_N_ON_OFF_2_O,
output   wire   [2:0]                                    out_N_ON_OFF_3_O,
//south ports														 
output   wire   [(3*flit_width)-1:0]                     out_S_FLIT_o,
output   wire   [2:0]                                    out_S_VALID_O,
output   wire   [2:0]                                    out_S_VC_0_RESERVED_O,
output   wire   [2:0]                                    out_S_VC_1_RESERVED_O,
output   wire   [2:0]                                    out_S_VC_2_RESERVED_O,
output   wire   [2:0]                                    out_S_VC_3_RESERVED_O,
output   wire   [2:0]                                    out_S_ON_OFF_0_O,
output   wire   [2:0]                                    out_S_ON_OFF_1_O,
output   wire   [2:0]                                    out_S_ON_OFF_2_O,
output   wire   [2:0]                                    out_S_ON_OFF_3_O,
//weast ports														 
output   wire   [(3*flit_width)-1:0]                     out_W_FLIT_o,
output   wire   [2:0]                                    out_W_VALID_O,
output   wire   [2:0]                                    out_W_VC_0_RESERVED_O,
output   wire   [2:0]                                    out_W_VC_1_RESERVED_O,
output   wire   [2:0]                                    out_W_VC_2_RESERVED_O,
output   wire   [2:0]                                    out_W_VC_3_RESERVED_O,
output   wire   [2:0]                                    out_W_ON_OFF_0_O,
output   wire   [2:0]                                    out_W_ON_OFF_1_O,
output   wire   [2:0]                                    out_W_ON_OFF_2_O,
output   wire   [2:0]                                    out_W_ON_OFF_3_O,
//east ports														 
output   wire   [(3*flit_width)-1:0]                     out_E_FLIT_o,
output   wire   [2:0]                                    out_E_VALID_O,
output   wire   [2:0]                                    out_E_VC_0_RESERVED_O,
output   wire   [2:0]                                    out_E_VC_1_RESERVED_O,
output   wire   [2:0]                                    out_E_VC_2_RESERVED_O,
output   wire   [2:0]                                    out_E_VC_3_RESERVED_O,
output   wire   [2:0]                                    out_E_ON_OFF_0_O,
output   wire   [2:0]                                    out_E_ON_OFF_1_O,
output   wire   [2:0]                                    out_E_ON_OFF_2_O,
output   wire   [2:0]                                    out_E_ON_OFF_3_O

);


///////////////////////instantiation////////////////////////////////////////

router_instanciate NOC_TOP (
.clk(clk),                  
.rst(rst),
.PE_VALID_i(PE_VALID_i),
.PE_FLIT_i(PE_FLIT_i),
.PE_VC_0_RESERVED_i(PE_VC_0_RESERVED_i),
.PE_VC_1_RESERVED_i(PE_VC_1_RESERVED_i),
.PE_VC_2_RESERVED_i(PE_VC_2_RESERVED_i),
.PE_VC_3_RESERVED_i(PE_VC_3_RESERVED_i),
.PE_ON_OFF_0_i(PE_ON_OFF_0_i),
.PE_ON_OFF_1_i(PE_ON_OFF_1_i),
.PE_ON_OFF_2_i(PE_ON_OFF_2_i),
.PE_ON_OFF_3_i(PE_ON_OFF_3_i),
.in_N_FLIT_i(in_N_FLIT_i),
.in_N_VALID_i(in_N_VALID_i),        
.in_N_VC_0_RESERVED_i(in_N_VC_0_RESERVED_i),
.in_N_VC_1_RESERVED_i(in_N_VC_1_RESERVED_i),
.in_N_VC_2_RESERVED_i(in_N_VC_2_RESERVED_i),
.in_N_VC_3_RESERVED_i(in_N_VC_3_RESERVED_i),
.in_N_ON_OFF_0_i(in_N_ON_OFF_0_i),
.in_N_ON_OFF_1_i(in_N_ON_OFF_1_i),
.in_N_ON_OFF_2_i(in_N_ON_OFF_2_i),
.in_N_ON_OFF_3_i(in_N_ON_OFF_3_i),
.in_S_FLIT_i(in_S_FLIT_i),
.in_S_VALID_i(in_S_VALID_i),        
.in_S_VC_0_RESERVED_i(in_S_VC_0_RESERVED_i),
.in_S_VC_1_RESERVED_i(in_S_VC_1_RESERVED_i),
.in_S_VC_2_RESERVED_i(in_S_VC_2_RESERVED_i),
.in_S_VC_3_RESERVED_i(in_S_VC_3_RESERVED_i),
.in_S_ON_OFF_0_i(in_S_ON_OFF_0_i),
.in_S_ON_OFF_1_i(in_S_ON_OFF_1_i),
.in_S_ON_OFF_2_i(in_S_ON_OFF_2_i),
.in_S_ON_OFF_3_i(in_S_ON_OFF_3_i),
.in_W_FLIT_i(in_W_FLIT_i),
.in_W_VALID_i(in_W_VALID_i),        
.in_W_VC_0_RESERVED_i(in_W_VC_0_RESERVED_i),
.in_W_VC_1_RESERVED_i(in_W_VC_1_RESERVED_i),
.in_W_VC_2_RESERVED_i(in_W_VC_2_RESERVED_i),
.in_W_VC_3_RESERVED_i(in_W_VC_3_RESERVED_i),
.in_W_ON_OFF_0_i(in_W_ON_OFF_0_i),
.in_W_ON_OFF_1_i(in_W_ON_OFF_1_i),
.in_W_ON_OFF_2_i(in_W_ON_OFF_2_i),
.in_W_ON_OFF_3_i(in_W_ON_OFF_3_i),
.in_E_FLIT_i(in_E_FLIT_i),
.in_E_VALID_i(in_E_VALID_i),        
.in_E_VC_0_RESERVED_i(in_E_VC_0_RESERVED_i),
.in_E_VC_1_RESERVED_i(in_E_VC_1_RESERVED_i),
.in_E_VC_2_RESERVED_i(in_E_VC_2_RESERVED_i),
.in_E_VC_3_RESERVED_i(in_E_VC_3_RESERVED_i),
.in_E_ON_OFF_0_i(in_E_ON_OFF_0_i),
.in_E_ON_OFF_1_i(in_E_ON_OFF_1_i),
.in_E_ON_OFF_2_i(in_E_ON_OFF_2_i),
.in_E_ON_OFF_3_i(in_E_ON_OFF_3_i),
.PE_FLIT_o(PE_FLIT_o),               
.PE_VALID_O(PE_VALID_O),
.PE_VC_0_RESERVED_O(PE_VC_0_RESERVED_O),
.PE_VC_1_RESERVED_O(PE_VC_1_RESERVED_O),
.PE_VC_2_RESERVED_O(PE_VC_2_RESERVED_O),
.PE_VC_3_RESERVED_O(PE_VC_3_RESERVED_O),
.PE_ON_OFF_0_O(PE_ON_OFF_0_O),
.PE_ON_OFF_1_O(PE_ON_OFF_1_O),
.PE_ON_OFF_2_O(PE_ON_OFF_2_O),
.PE_ON_OFF_3_O(PE_ON_OFF_3_O),
.out_N_FLIT_o(out_N_FLIT_o),
.out_N_VALID_O(out_N_VALID_O),
.out_N_VC_0_RESERVED_O(out_N_VC_0_RESERVED_O),
.out_N_VC_1_RESERVED_O(out_N_VC_1_RESERVED_O),
.out_N_VC_2_RESERVED_O(out_N_VC_2_RESERVED_O),
.out_N_VC_3_RESERVED_O(out_N_VC_3_RESERVED_O),
.out_N_ON_OFF_0_O(out_N_ON_OFF_0_O),
.out_N_ON_OFF_1_O(out_N_ON_OFF_1_O),
.out_N_ON_OFF_2_O(out_N_ON_OFF_2_O),
.out_N_ON_OFF_3_O(out_N_ON_OFF_3_O),
.out_S_FLIT_o(out_S_FLIT_o),
.out_S_VALID_O(out_S_VALID_O),
.out_S_VC_0_RESERVED_O(out_S_VC_0_RESERVED_O),
.out_S_VC_1_RESERVED_O(out_S_VC_1_RESERVED_O),
.out_S_VC_2_RESERVED_O(out_S_VC_2_RESERVED_O),
.out_S_VC_3_RESERVED_O(out_S_VC_3_RESERVED_O),
.out_S_ON_OFF_0_O(out_S_ON_OFF_0_O),
.out_S_ON_OFF_1_O(out_S_ON_OFF_1_O),
.out_S_ON_OFF_2_O(out_S_ON_OFF_2_O),
.out_S_ON_OFF_3_O(out_S_ON_OFF_3_O),
.out_W_FLIT_o(out_W_FLIT_o),
.out_W_VALID_O(out_W_VALID_O),
.out_W_VC_0_RESERVED_O(out_W_VC_0_RESERVED_O),
.out_W_VC_1_RESERVED_O(out_W_VC_1_RESERVED_O),
.out_W_VC_2_RESERVED_O(out_W_VC_2_RESERVED_O),
.out_W_VC_3_RESERVED_O(out_W_VC_3_RESERVED_O),
.out_W_ON_OFF_0_O(out_W_ON_OFF_0_O),
.out_W_ON_OFF_1_O(out_W_ON_OFF_1_O),
.out_W_ON_OFF_2_O(out_W_ON_OFF_2_O),
.out_W_ON_OFF_3_O(out_W_ON_OFF_3_O),
.out_E_FLIT_o(out_E_FLIT_o),
.out_E_VALID_O(out_E_VALID_O),
.out_E_VC_0_RESERVED_O(out_E_VC_0_RESERVED_O),
.out_E_VC_1_RESERVED_O(out_E_VC_1_RESERVED_O),
.out_E_VC_2_RESERVED_O(out_E_VC_2_RESERVED_O),
.out_E_VC_3_RESERVED_O(out_E_VC_3_RESERVED_O),
.out_E_ON_OFF_0_O(out_E_ON_OFF_0_O),
.out_E_ON_OFF_1_O(out_E_ON_OFF_1_O),
.out_E_ON_OFF_2_O(out_E_ON_OFF_2_O),
.out_E_ON_OFF_3_O(out_E_ON_OFF_3_O)
);

endmodule